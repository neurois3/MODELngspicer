trr.spice

.model DIODE1 D (
.include model.txt
+ )

V1  n01 0   dc 0 pulse(0 -3 10n 0.1n 0.1n 50n 100n 1)
V2  n04 0   dc 21.2
R1  n01 n02 50
R2  n02 0   50
R3  n03 n04 2k
R4  n05 0   50
C1  n02 n03 0.01u
D1  n03 n05 DIODE1

.control
tran 10p 20n
wrdata trr.txt v(n05)
.endc
.end
