if-vf.spice

.model DIODE1 D (
.include model.txt
+ )

V1  n01 0   dc 0
D1  n01 0   DIODE1

.control
option TEMP=25
dc V1 0.3 1.5 0.01

set wr_singlescale
wrdata if-vf.txt -i(V1)
.endc
.end
