NMOS_ID_VDS.spice
* This script performs a DC sweep of VDS for multiple VGS values
* to extract the drain current (I_D) characteristics of an NMOS transistor.

.model NMOS1 NMOS (
+ level=1 L=1u W=100u
.include model.txt
+ )

* Voltage sources
VGS g   0           dc 0    $ Gate-to-Source voltage source
VDS dd  0           dc 0    $ Drain-to-Source voltage source
VID dd  d           dc 0    $ Current probe for I_D

* NMOS transistor instance
M1  d   g   0   0   NMOS1   $ Test NMOS transistor

.control
option TEMP=25              $ Set simulation temperature to 25°C
foreach VGS_value 1.4 1.5 1.7 1.9 2.0 2.5
    alter VGS dc = $VGS_value       $ Set VGS to current value
    dc VDS 0.1 15 0.01              $ Sweep VDS from 0.1 V to 15 V in 0.1 V steps
end

* Write drain current results to file
set wr_singlescale
wrdata NMOS_ID_VDS.txt
+ dc1.i(VID) dc2.i(VID) dc3.i(VID) dc4.i(VID)
+ dc5.i(VID) dc6.i(VID)  $ Drain current for each VGS sweep

.endc
.end
