ir-vr.spice

.model DIODE1 D (
.include model.txt
+ )

V1  n01 0   dc 0
D1  0   n01 DIODE1

.control
option TEMP=25 GMIN=4e-10
dc V1 10 146 1

set wr_singlescale
wrdata ir-vr.txt -i(V1)
.endc
.end
