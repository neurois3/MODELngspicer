NMOS_ID_VGS.spice
* This script performs a DC sweep of VGS at a fixed VDS
* to extract the drain current (I_D) vs. gate voltage characteristics.

.model NMOS1 NMOS (
+ level=1 L=1u W=100u
.include model.txt
+ )

* Voltage sources
VGS g   0           dc 0    $ Gate-to-Source voltage source
VDS dd  0           dc 15   $ Drain-to-Source voltage source
VID dd  d           dc 0    $ Current probe for I_D

* NMOS transistor instance
M1  d   g   0   0   NMOS1   $ Test NMOS transistor

.control
option TEMP=25              $ Set simulation temperature to 25°C

* Sweep VGS from 1.3 V to 2.5 V in 0.01 V steps
dc VGS 1.3 2.5 0.01

* Write drain current results to file
set wr_singlescale
wrdata NMOS_ID_VGS.txt i(VID)

.endc
.end
